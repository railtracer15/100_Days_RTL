`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Create Date: 18.03.2025 09:50:08
// Module Name: N_bit_comp_tb
//////////////////////////////////////////////////////////////////////////////////


module N_bit_comp_tb(

    );
    parameter N=8;
    reg [N-1:0] A ,B ;
    wire gt ,ls ,eq ;
    N_bit_comp dut(.A(A),.B(B),.gt(gt),.ls(ls),.eq(eq));
    initial begin
        A = 8'b10100001; B = 8'b10100001;
        #10;
        A = 8'b00001100; B = 8'b00001010;
        #10;
        A = 8'b00000011; B = 8'b00000100;
        #10;
        A = 8'b00000000; B = 8'b00000000;
        #10;
        A = 8'b11111111; B = 8'b01111111;
        #10;
        A = 8'b00000001; B = 8'b00000010;
        #10;
        $finish;
    end
    
endmodule
